class scoreboard extends uvm_scoreboard;
  `uvm_component_utils(scoreboard)
    
endclass
 
